// Description
`timescale 1ns / 1ps

module project_LED_blink_tb();

endmodule